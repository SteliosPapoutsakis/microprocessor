module Data_path(Addr_out,Addr_in,Valid,regEn,oppB,oppA,opcode,fetch,literal)

endmodule //
