package common;
typedef enum {S_fetch,S_Decode,S_ExecuteArth,S_ExecuteLS,S_ExecuteBR,S_store} motherStates;
typedef enum {State1,State2,State3,State4,State5,State6,State7,State8,State9} States;
endpackage
